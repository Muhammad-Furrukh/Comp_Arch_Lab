import cep_define ::*;
module addr_check_n_tb();
  logic unsigned [31:0]addr, addr_n,addr_n_1;
  logic [1:0]size;
  logic [1:0] a_n;
  logic out;

  addr_check_n DUT(.*);

  initial begin
    // Testing for OFF mode
    addr_n = 32'h1234567E; addr_n_1 = 32'h1234566E; addr = 32'h1234566D; size = 2'b00; a_n = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h1234566E; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h1234567D; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h1234567E; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;

    // Testing for TOR mode
    addr = 32'h1234566D; size = 2'b00; a_n = 2'b01;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h1234566E; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h1234567D; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h1234567E; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;

    // Testing for NA4 mode
    addr = 32'h1234566D; size = 2'b00; a_n = 2'b10;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h1234566E; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h1234567D; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h1234567E; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h1234567F; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h12345680; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h12345681; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = 32'h12345682; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;

    // Testing for NAPOT mode
    addr = (32'h1234566E & (~(32'b1))) - 1; size = 2'b00; a_n = 2'b11;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = (32'h1234566E & (~(32'b1))); size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = (32'h1234567E & (~(32'b1))) - 1; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = (32'h1234567E & (~(32'b1))); size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = (32'h1234567E & (~(32'b1))) + 7; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    addr = (32'h1234567E & (~(32'b1))) + 8; size = 2'b00;
    #10;
    size = 2'b01;
    #10;
    size = 2'b11;
    #10;
    $stop;
  end
endmodule