module Tx_Cont_Stat_Reg();

endmodule