module UART_Tx_tb();

endmodule